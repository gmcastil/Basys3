module user_core //#(
//)
(
);

endmodule

